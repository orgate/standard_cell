magic
tech sample_6m
timestamp 1384533072
<< nwell >>
rect -11 32 61 76
<< pwell >>
rect -11 -4 61 32
<< ntransistor >>
rect 6 15 8 25
rect 15 15 17 25
rect 24 15 26 25
rect 33 15 35 24
<< ptransistor >>
rect 6 38 8 58
rect 15 38 17 58
rect 24 38 26 58
rect 33 38 35 58
rect 42 38 44 48
<< ndiffusion >>
rect 5 15 6 25
rect 8 15 9 25
rect 14 15 15 25
rect 17 15 18 25
rect 23 15 24 25
rect 26 15 27 25
rect 32 15 33 24
rect 35 15 36 24
<< pdiffusion >>
rect 5 38 6 58
rect 8 38 9 58
rect 14 38 15 58
rect 17 38 18 58
rect 23 38 24 58
rect 26 38 27 58
rect 32 38 33 58
rect 35 38 36 58
rect 41 38 42 48
rect 44 38 45 48
<< ndcontact >>
rect 0 15 5 25
rect 9 15 14 25
rect 18 15 23 25
rect 27 15 32 25
rect 36 15 41 24
<< pdcontact >>
rect 0 38 5 58
rect 9 38 14 58
rect 18 38 23 58
rect 27 38 32 58
rect 36 38 41 58
rect 45 38 50 48
<< psubstratepcontact >>
rect 52 1 60 7
<< nsubstratencontact >>
rect 52 65 60 71
<< polysilicon >>
rect 6 58 8 61
rect 15 58 17 61
rect 24 58 26 61
rect 33 58 35 61
rect 42 48 44 51
rect 6 36 8 38
rect 15 36 17 38
rect 24 36 26 38
rect 33 36 35 38
rect 42 36 44 38
rect 6 34 44 36
rect -1 30 2 34
rect 6 25 8 34
rect 15 25 17 34
rect 24 25 26 34
rect 33 24 35 34
rect 6 12 8 15
rect 15 12 17 15
rect 24 12 26 15
rect 33 12 35 15
rect 42 12 44 34
<< polycontact >>
rect -5 30 -1 34
rect 2 30 6 34
<< metal1 >>
rect -11 64 61 72
rect 0 58 5 64
rect 18 58 23 64
rect 36 58 41 64
rect -9 30 -5 34
rect 9 31 14 38
rect 27 31 32 38
rect 45 31 50 38
rect 9 28 50 31
rect 9 25 14 28
rect 27 25 32 28
rect 0 8 5 15
rect 18 8 23 15
rect 36 8 41 15
rect -11 7 61 8
rect -11 1 52 7
rect 60 1 61 7
rect -11 0 61 1
<< labels >>
rlabel metal1 19 69 22 72 5 Vdd 
rlabel metal1 19 0 21 3 1 Gnd
rlabel metal1 -9 31 -8 32 3 in
rlabel metal1 13 29 14 30 1 out
<< end >>
